library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

use work.StatePackage.all;

entity VGA40 is
    Port ( clock_50      : in  STD_LOGIC;
           reset         : in  STD_LOGIC;
           Hsync         : out STD_LOGIC;
           Vsync         : out STD_LOGIC;
           vga_r         : out STD_LOGIC_VECTOR (11 downto 0);
           vga_g         : out STD_LOGIC_VECTOR (11 downto 0);
           vga_b         : out STD_LOGIC_VECTOR (11 downto 0);
           vga_hs        : out STD_LOGIC;
           vga_vs        : out STD_LOGIC;
			  current_state : in state 
			 );
end VGA40;

architecture Behavioral of VGA40 is

-- VGA Controller constants
constant HOR_RES    : integer := 640;   -- Horizontal resolution
constant VER_RES    : integer := 480;   -- Vertical resolution
constant HOR_FRONT  : integer := 16;    -- Horizontal Front Porch
constant HOR_SYNC   : integer := 96;    -- Horizontal Sync pulse width
constant HOR_BACK   : integer := 48;    -- Horizontal Back Porch
constant VER_FRONT  : integer := 10;    -- Vertical Front Porch
constant VER_SYNC   : integer := 2;     -- Vertical Sync pulse width
constant VER_BACK   : integer := 33;    -- Vertical Back Porch

-- 12-bit Sine LUT
type SIN_LUT_TYPE is array (0 to 4095) of STD_LOGIC_VECTOR(11 downto 0);
constant SIN_LUT : SIN_LUT_TYPE := (
"011111111111","100000000010","100000000101","100000001000","100000001100","100000001111","100000010010","100000010101",
"100000011000","100000011011","100000011110","100000100010","100000100101","100000101000","100000101011","100000101110",
"100000110001","100000110100","100000111000","100000111011","100000111110","100001000001","100001000100","100001000111",
"100001001010","100001001110","100001010001","100001010100","100001010111","100001011010","100001011101","100001100000",
"100001100011","100001100111","100001101010","100001101101","100001110000","100001110011","100001110110","100001111001",
"100001111101","100010000000","100010000011","100010000110","100010001001","100010001100","100010001111","100010010010",
"100010010110","100010011001","100010011100","100010011111","100010100010","100010100101","100010101000","100010101100",
"100010101111","100010110010","100010110101","100010111000","100010111011","100010111110","100011000001","100011000101",
"100011001000","100011001011","100011001110","100011010001","100011010100","100011010111","100011011010","100011011110",
"100011100001","100011100100","100011100111","100011101010","100011101101","100011110000","100011110011","100011110111",
"100011111010","100011111101","100100000000","100100000011","100100000110","100100001001","100100001100","100100001111",
"100100010011","100100010110","100100011001","100100011100","100100011111","100100100010","100100100101","100100101000",
"100100101011","100100101111","100100110010","100100110101","100100111000","100100111011","100100111110","100101000001",
"100101000100","100101000111","100101001010","100101001110","100101010001","100101010100","100101010111","100101011010",
"100101011101","100101100000","100101100011","100101100110","100101101001","100101101101","100101110000","100101110011",
"100101110110","100101111001","100101111100","100101111111","100110000010","100110000101","100110001000","100110001011",
"100110001110","100110010010","100110010101","100110011000","100110011011","100110011110","100110100001","100110100100",
"100110100111","100110101010","100110101101","100110110000","100110110011","100110110110","100110111001","100110111101",
"100111000000","100111000011","100111000110","100111001001","100111001100","100111001111","100111010010","100111010101",
"100111011000","100111011011","100111011110","100111100001","100111100100","100111100111","100111101010","100111101101",
"100111110001","100111110100","100111110111","100111111010","100111111101","101000000000","101000000011","101000000110",
"101000001001","101000001100","101000001111","101000010010","101000010101","101000011000","101000011011","101000011110",
"101000100001","101000100100","101000100111","101000101010","101000101101","101000110000","101000110011","101000110110",
"101000111001","101000111100","101000111111","101001000010","101001000101","101001001000","101001001011","101001001110",
"101001010001","101001010100","101001010111","101001011010","101001011101","101001100000","101001100011","101001100110",
"101001101001","101001101100","101001101111","101001110010","101001110101","101001111000","101001111011","101001111110",
"101010000001","101010000100","101010000111","101010001010","101010001101","101010010000","101010010011","101010010110",
"101010011001","101010011100","101010011111","101010100010","101010100101","101010101000","101010101011","101010101110",
"101010110001","101010110100","101010110111","101010111010","101010111101","101011000000","101011000010","101011000101",
"101011001000","101011001011","101011001110","101011010001","101011010100","101011010111","101011011010","101011011101",
"101011100000","101011100011","101011100110","101011101001","101011101100","101011101111","101011110001","101011110100",
"101011110111","101011111010","101011111101","101100000000","101100000011","101100000110","101100001001","101100001100",
"101100001111","101100010001","101100010100","101100010111","101100011010","101100011101","101100100000","101100100011",
"101100100110","101100101001","101100101011","101100101110","101100110001","101100110100","101100110111","101100111010",
"101100111101","101101000000","101101000010","101101000101","101101001000","101101001011","101101001110","101101010001",
"101101010100","101101010110","101101011001","101101011100","101101011111","101101100010","101101100101","101101101000",
"101101101010","101101101101","101101110000","101101110011","101101110110","101101111001","101101111011","101101111110",
"101110000001","101110000100","101110000111","101110001010","101110001100","101110001111","101110010010","101110010101",
"101110011000","101110011010","101110011101","101110100000","101110100011","101110100110","101110101000","101110101011",
"101110101110","101110110001","101110110100","101110110110","101110111001","101110111100","101110111111","101111000001",
"101111000100","101111000111","101111001010","101111001100","101111001111","101111010010","101111010101","101111011000",
"101111011010","101111011101","101111100000","101111100011","101111100101","101111101000","101111101011","101111101101",
"101111110000","101111110011","101111110110","101111111000","101111111011","101111111110","110000000001","110000000011",
"110000000110","110000001001","110000001011","110000001110","110000010001","110000010100","110000010110","110000011001",
"110000011100","110000011110","110000100001","110000100100","110000100110","110000101001","110000101100","110000101110",
"110000110001","110000110100","110000110110","110000111001","110000111100","110000111110","110001000001","110001000100",
"110001000110","110001001001","110001001100","110001001110","110001010001","110001010100","110001010110","110001011001",
"110001011100","110001011110","110001100001","110001100011","110001100110","110001101001","110001101011","110001101110",
"110001110001","110001110011","110001110110","110001111000","110001111011","110001111110","110010000000","110010000011",
"110010000101","110010001000","110010001011","110010001101","110010010000","110010010010","110010010101","110010010111",
"110010011010","110010011101","110010011111","110010100010","110010100100","110010100111","110010101001","110010101100",
"110010101110","110010110001","110010110100","110010110110","110010111001","110010111011","110010111110","110011000000",
"110011000011","110011000101","110011001000","110011001010","110011001101","110011001111","110011010010","110011010100",
"110011010111","110011011001","110011011100","110011011110","110011100001","110011100011","110011100110","110011101000",
"110011101011","110011101101","110011110000","110011110010","110011110101","110011110111","110011111001","110011111100",
"110011111110","110100000001","110100000011","110100000110","110100001000","110100001011","110100001101","110100001111",
"110100010010","110100010100","110100010111","110100011001","110100011100","110100011110","110100100000","110100100011",
"110100100101","110100101000","110100101010","110100101100","110100101111","110100110001","110100110100","110100110110",
"110100111000","110100111011","110100111101","110100111111","110101000010","110101000100","110101000111","110101001001",
"110101001011","110101001110","110101010000","110101010010","110101010101","110101010111","110101011001","110101011100",
"110101011110","110101100000","110101100011","110101100101","110101100111","110101101010","110101101100","110101101110",
"110101110001","110101110011","110101110101","110101110111","110101111010","110101111100","110101111110","110110000001",
"110110000011","110110000101","110110000111","110110001010","110110001100","110110001110","110110010000","110110010011",
"110110010101","110110010111","110110011001","110110011100","110110011110","110110100000","110110100010","110110100101",
"110110100111","110110101001","110110101011","110110101101","110110110000","110110110010","110110110100","110110110110",
"110110111000","110110111011","110110111101","110110111111","110111000001","110111000011","110111000110","110111001000",
"110111001010","110111001100","110111001110","110111010000","110111010011","110111010101","110111010111","110111011001",
"110111011011","110111011101","110111011111","110111100010","110111100100","110111100110","110111101000","110111101010",
"110111101100","110111101110","110111110000","110111110010","110111110101","110111110111","110111111001","110111111011",
"110111111101","110111111111","111000000001","111000000011","111000000101","111000000111","111000001001","111000001011",
"111000001101","111000001111","111000010001","111000010100","111000010110","111000011000","111000011010","111000011100",
"111000011110","111000100000","111000100010","111000100100","111000100110","111000101000","111000101010","111000101100",
"111000101110","111000110000","111000110010","111000110100","111000110110","111000111000","111000111010","111000111100",
"111000111110","111001000000","111001000001","111001000011","111001000101","111001000111","111001001001","111001001011",
"111001001101","111001001111","111001010001","111001010011","111001010101","111001010111","111001011001","111001011011",
"111001011100","111001011110","111001100000","111001100010","111001100100","111001100110","111001101000","111001101010",
"111001101100","111001101101","111001101111","111001110001","111001110011","111001110101","111001110111","111001111001",
"111001111010","111001111100","111001111110","111010000000","111010000010","111010000100","111010000101","111010000111",
"111010001001","111010001011","111010001101","111010001110","111010010000","111010010010","111010010100","111010010110",
"111010010111","111010011001","111010011011","111010011101","111010011110","111010100000","111010100010","111010100100",
"111010100101","111010100111","111010101001","111010101011","111010101100","111010101110","111010110000","111010110010",
"111010110011","111010110101","111010110111","111010111000","111010111010","111010111100","111010111101","111010111111",
"111011000001","111011000011","111011000100","111011000110","111011001000","111011001001","111011001011","111011001101",
"111011001110","111011010000","111011010001","111011010011","111011010101","111011010110","111011011000","111011011010",
"111011011011","111011011101","111011011110","111011100000","111011100010","111011100011","111011100101","111011100110",
"111011101000","111011101010","111011101011","111011101101","111011101110","111011110000","111011110001","111011110011",
"111011110101","111011110110","111011111000","111011111001","111011111011","111011111100","111011111110","111011111111",
"111100000001","111100000010","111100000100","111100000101","111100000111","111100001000","111100001010","111100001011",
"111100001101","111100001110","111100010000","111100010001","111100010011","111100010100","111100010110","111100010111",
"111100011000","111100011010","111100011011","111100011101","111100011110","111100100000","111100100001","111100100010",
"111100100100","111100100101","111100100111","111100101000","111100101001","111100101011","111100101100","111100101110",
"111100101111","111100110000","111100110010","111100110011","111100110101","111100110110","111100110111","111100111001",
"111100111010","111100111011","111100111101","111100111110","111100111111","111101000001","111101000010","111101000011",
"111101000101","111101000110","111101000111","111101001000","111101001010","111101001011","111101001100","111101001110",
"111101001111","111101010000","111101010001","111101010011","111101010100","111101010101","111101010110","111101011000",
"111101011001","111101011010","111101011011","111101011101","111101011110","111101011111","111101100000","111101100001",
"111101100011","111101100100","111101100101","111101100110","111101100111","111101101001","111101101010","111101101011",
"111101101100","111101101101","111101101110","111101110000","111101110001","111101110010","111101110011","111101110100",
"111101110101","111101110110","111101111000","111101111001","111101111010","111101111011","111101111100","111101111101",
"111101111110","111101111111","111110000000","111110000001","111110000011","111110000100","111110000101","111110000110",
"111110000111","111110001000","111110001001","111110001010","111110001011","111110001100","111110001101","111110001110",
"111110001111","111110010000","111110010001","111110010010","111110010011","111110010100","111110010101","111110010110",
"111110010111","111110011000","111110011001","111110011010","111110011011","111110011100","111110011101","111110011110",
"111110011111","111110100000","111110100001","111110100010","111110100011","111110100100","111110100101","111110100101",
"111110100110","111110100111","111110101000","111110101001","111110101010","111110101011","111110101100","111110101101",
"111110101101","111110101110","111110101111","111110110000","111110110001","111110110010","111110110011","111110110011",
"111110110100","111110110101","111110110110","111110110111","111110111000","111110111000","111110111001","111110111010",
"111110111011","111110111100","111110111100","111110111101","111110111110","111110111111","111111000000","111111000000",
"111111000001","111111000010","111111000011","111111000011","111111000100","111111000101","111111000110","111111000110",
"111111000111","111111001000","111111001001","111111001001","111111001010","111111001011","111111001011","111111001100",
"111111001101","111111001101","111111001110","111111001111","111111001111","111111010000","111111010001","111111010001",
"111111010010","111111010011","111111010011","111111010100","111111010101","111111010101","111111010110","111111010111",
"111111010111","111111011000","111111011000","111111011001","111111011010","111111011010","111111011011","111111011011",
"111111011100","111111011100","111111011101","111111011110","111111011110","111111011111","111111011111","111111100000",
"111111100000","111111100001","111111100001","111111100010","111111100010","111111100011","111111100011","111111100100",
"111111100100","111111100101","111111100101","111111100110","111111100110","111111100111","111111100111","111111101000",
"111111101000","111111101001","111111101001","111111101010","111111101010","111111101011","111111101011","111111101011",
"111111101100","111111101100","111111101101","111111101101","111111101110","111111101110","111111101110","111111101111",
"111111101111","111111101111","111111110000","111111110000","111111110001","111111110001","111111110001","111111110010",
"111111110010","111111110010","111111110011","111111110011","111111110011","111111110100","111111110100","111111110100",
"111111110101","111111110101","111111110101","111111110110","111111110110","111111110110","111111110110","111111110111",
"111111110111","111111110111","111111110111","111111111000","111111111000","111111111000","111111111000","111111111001",
"111111111001","111111111001","111111111001","111111111010","111111111010","111111111010","111111111010","111111111010",
"111111111011","111111111011","111111111011","111111111011","111111111011","111111111100","111111111100","111111111100",
"111111111100","111111111100","111111111100","111111111100","111111111101","111111111101","111111111101","111111111101",
"111111111101","111111111101","111111111101","111111111101","111111111110","111111111110","111111111110","111111111110",
"111111111110","111111111110","111111111110","111111111110","111111111110","111111111110","111111111110","111111111110",
"111111111110","111111111110","111111111110","111111111110","111111111110","111111111110","111111111110","111111111110",
"111111111111","111111111110","111111111110","111111111110","111111111110","111111111110","111111111110","111111111110",
"111111111110","111111111110","111111111110","111111111110","111111111110","111111111110","111111111110","111111111110",
"111111111110","111111111110","111111111110","111111111110","111111111110","111111111101","111111111101","111111111101",
"111111111101","111111111101","111111111101","111111111101","111111111101","111111111100","111111111100","111111111100",
"111111111100","111111111100","111111111100","111111111100","111111111011","111111111011","111111111011","111111111011",
"111111111011","111111111010","111111111010","111111111010","111111111010","111111111010","111111111001","111111111001",
"111111111001","111111111001","111111111000","111111111000","111111111000","111111111000","111111110111","111111110111",
"111111110111","111111110111","111111110110","111111110110","111111110110","111111110110","111111110101","111111110101",
"111111110101","111111110100","111111110100","111111110100","111111110011","111111110011","111111110011","111111110010",
"111111110010","111111110010","111111110001","111111110001","111111110001","111111110000","111111110000","111111101111",
"111111101111","111111101111","111111101110","111111101110","111111101110","111111101101","111111101101","111111101100",
"111111101100","111111101011","111111101011","111111101011","111111101010","111111101010","111111101001","111111101001",
"111111101000","111111101000","111111100111","111111100111","111111100110","111111100110","111111100101","111111100101",
"111111100100","111111100100","111111100011","111111100011","111111100010","111111100010","111111100001","111111100001",
"111111100000","111111100000","111111011111","111111011111","111111011110","111111011110","111111011101","111111011100",
"111111011100","111111011011","111111011011","111111011010","111111011010","111111011001","111111011000","111111011000",
"111111010111","111111010111","111111010110","111111010101","111111010101","111111010100","111111010011","111111010011",
"111111010010","111111010001","111111010001","111111010000","111111001111","111111001111","111111001110","111111001101",
"111111001101","111111001100","111111001011","111111001011","111111001010","111111001001","111111001001","111111001000",
"111111000111","111111000110","111111000110","111111000101","111111000100","111111000011","111111000011","111111000010",
"111111000001","111111000000","111111000000","111110111111","111110111110","111110111101","111110111100","111110111100",
"111110111011","111110111010","111110111001","111110111000","111110111000","111110110111","111110110110","111110110101",
"111110110100","111110110011","111110110011","111110110010","111110110001","111110110000","111110101111","111110101110",
"111110101101","111110101101","111110101100","111110101011","111110101010","111110101001","111110101000","111110100111",
"111110100110","111110100101","111110100101","111110100100","111110100011","111110100010","111110100001","111110100000",
"111110011111","111110011110","111110011101","111110011100","111110011011","111110011010","111110011001","111110011000",
"111110010111","111110010110","111110010101","111110010100","111110010011","111110010010","111110010001","111110010000",
"111110001111","111110001110","111110001101","111110001100","111110001011","111110001010","111110001001","111110001000",
"111110000111","111110000110","111110000101","111110000100","111110000011","111110000001","111110000000","111101111111",
"111101111110","111101111101","111101111100","111101111011","111101111010","111101111001","111101111000","111101110110",
"111101110101","111101110100","111101110011","111101110010","111101110001","111101110000","111101101110","111101101101",
"111101101100","111101101011","111101101010","111101101001","111101100111","111101100110","111101100101","111101100100",
"111101100011","111101100001","111101100000","111101011111","111101011110","111101011101","111101011011","111101011010",
"111101011001","111101011000","111101010110","111101010101","111101010100","111101010011","111101010001","111101010000",
"111101001111","111101001110","111101001100","111101001011","111101001010","111101001000","111101000111","111101000110",
"111101000101","111101000011","111101000010","111101000001","111100111111","111100111110","111100111101","111100111011",
"111100111010","111100111001","111100110111","111100110110","111100110101","111100110011","111100110010","111100110000",
"111100101111","111100101110","111100101100","111100101011","111100101001","111100101000","111100100111","111100100101",
"111100100100","111100100010","111100100001","111100100000","111100011110","111100011101","111100011011","111100011010",
"111100011000","111100010111","111100010110","111100010100","111100010011","111100010001","111100010000","111100001110",
"111100001101","111100001011","111100001010","111100001000","111100000111","111100000101","111100000100","111100000010",
"111100000001","111011111111","111011111110","111011111100","111011111011","111011111001","111011111000","111011110110",
"111011110101","111011110011","111011110001","111011110000","111011101110","111011101101","111011101011","111011101010",
"111011101000","111011100110","111011100101","111011100011","111011100010","111011100000","111011011110","111011011101",
"111011011011","111011011010","111011011000","111011010110","111011010101","111011010011","111011010001","111011010000",
"111011001110","111011001101","111011001011","111011001001","111011001000","111011000110","111011000100","111011000011",
"111011000001","111010111111","111010111101","111010111100","111010111010","111010111000","111010110111","111010110101",
"111010110011","111010110010","111010110000","111010101110","111010101100","111010101011","111010101001","111010100111",
"111010100101","111010100100","111010100010","111010100000","111010011110","111010011101","111010011011","111010011001",
"111010010111","111010010110","111010010100","111010010010","111010010000","111010001110","111010001101","111010001011",
"111010001001","111010000111","111010000101","111010000100","111010000010","111010000000","111001111110","111001111100",
"111001111010","111001111001","111001110111","111001110101","111001110011","111001110001","111001101111","111001101101",
"111001101100","111001101010","111001101000","111001100110","111001100100","111001100010","111001100000","111001011110",
"111001011100","111001011011","111001011001","111001010111","111001010101","111001010011","111001010001","111001001111",
"111001001101","111001001011","111001001001","111001000111","111001000101","111001000011","111001000001","111001000000",
"111000111110","111000111100","111000111010","111000111000","111000110110","111000110100","111000110010","111000110000",
"111000101110","111000101100","111000101010","111000101000","111000100110","111000100100","111000100010","111000100000",
"111000011110","111000011100","111000011010","111000011000","111000010110","111000010100","111000010001","111000001111",
"111000001101","111000001011","111000001001","111000000111","111000000101","111000000011","111000000001","110111111111",
"110111111101","110111111011","110111111001","110111110111","110111110101","110111110010","110111110000","110111101110",
"110111101100","110111101010","110111101000","110111100110","110111100100","110111100010","110111011111","110111011101",
"110111011011","110111011001","110111010111","110111010101","110111010011","110111010000","110111001110","110111001100",
"110111001010","110111001000","110111000110","110111000011","110111000001","110110111111","110110111101","110110111011",
"110110111000","110110110110","110110110100","110110110010","110110110000","110110101101","110110101011","110110101001",
"110110100111","110110100101","110110100010","110110100000","110110011110","110110011100","110110011001","110110010111",
"110110010101","110110010011","110110010000","110110001110","110110001100","110110001010","110110000111","110110000101",
"110110000011","110110000001","110101111110","110101111100","110101111010","110101110111","110101110101","110101110011",
"110101110001","110101101110","110101101100","110101101010","110101100111","110101100101","110101100011","110101100000",
"110101011110","110101011100","110101011001","110101010111","110101010101","110101010010","110101010000","110101001110",
"110101001011","110101001001","110101000111","110101000100","110101000010","110100111111","110100111101","110100111011",
"110100111000","110100110110","110100110100","110100110001","110100101111","110100101100","110100101010","110100101000",
"110100100101","110100100011","110100100000","110100011110","110100011100","110100011001","110100010111","110100010100",
"110100010010","110100001111","110100001101","110100001011","110100001000","110100000110","110100000011","110100000001",
"110011111110","110011111100","110011111001","110011110111","110011110101","110011110010","110011110000","110011101101",
"110011101011","110011101000","110011100110","110011100011","110011100001","110011011110","110011011100","110011011001",
"110011010111","110011010100","110011010010","110011001111","110011001101","110011001010","110011001000","110011000101",
"110011000011","110011000000","110010111110","110010111011","110010111001","110010110110","110010110100","110010110001",
"110010101110","110010101100","110010101001","110010100111","110010100100","110010100010","110010011111","110010011101",
"110010011010","110010010111","110010010101","110010010010","110010010000","110010001101","110010001011","110010001000",
"110010000101","110010000011","110010000000","110001111110","110001111011","110001111000","110001110110","110001110011",
"110001110001","110001101110","110001101011","110001101001","110001100110","110001100011","110001100001","110001011110",
"110001011100","110001011001","110001010110","110001010100","110001010001","110001001110","110001001100","110001001001",
"110001000110","110001000100","110001000001","110000111110","110000111100","110000111001","110000110110","110000110100",
"110000110001","110000101110","110000101100","110000101001","110000100110","110000100100","110000100001","110000011110",
"110000011100","110000011001","110000010110","110000010100","110000010001","110000001110","110000001011","110000001001",
"110000000110","110000000011","110000000001","101111111110","101111111011","101111111000","101111110110","101111110011",
"101111110000","101111101101","101111101011","101111101000","101111100101","101111100011","101111100000","101111011101",
"101111011010","101111011000","101111010101","101111010010","101111001111","101111001100","101111001010","101111000111",
"101111000100","101111000001","101110111111","101110111100","101110111001","101110110110","101110110100","101110110001",
"101110101110","101110101011","101110101000","101110100110","101110100011","101110100000","101110011101","101110011010",
"101110011000","101110010101","101110010010","101110001111","101110001100","101110001010","101110000111","101110000100",
"101110000001","101101111110","101101111011","101101111001","101101110110","101101110011","101101110000","101101101101",
"101101101010","101101101000","101101100101","101101100010","101101011111","101101011100","101101011001","101101010110",
"101101010100","101101010001","101101001110","101101001011","101101001000","101101000101","101101000010","101101000000",
"101100111101","101100111010","101100110111","101100110100","101100110001","101100101110","101100101011","101100101001",
"101100100110","101100100011","101100100000","101100011101","101100011010","101100010111","101100010100","101100010001",
"101100001111","101100001100","101100001001","101100000110","101100000011","101100000000","101011111101","101011111010",
"101011110111","101011110100","101011110001","101011101111","101011101100","101011101001","101011100110","101011100011",
"101011100000","101011011101","101011011010","101011010111","101011010100","101011010001","101011001110","101011001011",
"101011001000","101011000101","101011000010","101011000000","101010111101","101010111010","101010110111","101010110100",
"101010110001","101010101110","101010101011","101010101000","101010100101","101010100010","101010011111","101010011100",
"101010011001","101010010110","101010010011","101010010000","101010001101","101010001010","101010000111","101010000100",
"101010000001","101001111110","101001111011","101001111000","101001110101","101001110010","101001101111","101001101100",
"101001101001","101001100110","101001100011","101001100000","101001011101","101001011010","101001010111","101001010100",
"101001010001","101001001110","101001001011","101001001000","101001000101","101001000010","101000111111","101000111100",
"101000111001","101000110110","101000110011","101000110000","101000101101","101000101010","101000100111","101000100100",
"101000100001","101000011110","101000011011","101000011000","101000010101","101000010010","101000001111","101000001100",
"101000001001","101000000110","101000000011","101000000000","100111111101","100111111010","100111110111","100111110100",
"100111110001","100111101101","100111101010","100111100111","100111100100","100111100001","100111011110","100111011011",
"100111011000","100111010101","100111010010","100111001111","100111001100","100111001001","100111000110","100111000011",
"100111000000","100110111101","100110111001","100110110110","100110110011","100110110000","100110101101","100110101010",
"100110100111","100110100100","100110100001","100110011110","100110011011","100110011000","100110010101","100110010010",
"100110001110","100110001011","100110001000","100110000101","100110000010","100101111111","100101111100","100101111001",
"100101110110","100101110011","100101110000","100101101101","100101101001","100101100110","100101100011","100101100000",
"100101011101","100101011010","100101010111","100101010100","100101010001","100101001110","100101001010","100101000111",
"100101000100","100101000001","100100111110","100100111011","100100111000","100100110101","100100110010","100100101111",
"100100101011","100100101000","100100100101","100100100010","100100011111","100100011100","100100011001","100100010110",
"100100010011","100100001111","100100001100","100100001001","100100000110","100100000011","100100000000","100011111101",
"100011111010","100011110111","100011110011","100011110000","100011101101","100011101010","100011100111","100011100100",
"100011100001","100011011110","100011011010","100011010111","100011010100","100011010001","100011001110","100011001011",
"100011001000","100011000101","100011000001","100010111110","100010111011","100010111000","100010110101","100010110010",
"100010101111","100010101100","100010101000","100010100101","100010100010","100010011111","100010011100","100010011001",
"100010010110","100010010010","100010001111","100010001100","100010001001","100010000110","100010000011","100010000000",
"100001111101","100001111001","100001110110","100001110011","100001110000","100001101101","100001101010","100001100111",
"100001100011","100001100000","100001011101","100001011010","100001010111","100001010100","100001010001","100001001110",
"100001001010","100001000111","100001000100","100001000001","100000111110","100000111011","100000111000","100000110100",
"100000110001","100000101110","100000101011","100000101000","100000100101","100000100010","100000011110","100000011011",
"100000011000","100000010101","100000010010","100000001111","100000001100","100000001000","100000000101","100000000010",
"011111111111","011111111100","011111111001","011111110110","011111110010","011111101111","011111101100","011111101001",
"011111100110","011111100011","011111100000","011111011100","011111011001","011111010110","011111010011","011111010000",
"011111001101","011111001010","011111000110","011111000011","011111000000","011110111101","011110111010","011110110111",
"011110110100","011110110000","011110101101","011110101010","011110100111","011110100100","011110100001","011110011110",
"011110011011","011110010111","011110010100","011110010001","011110001110","011110001011","011110001000","011110000101",
"011110000001","011101111110","011101111011","011101111000","011101110101","011101110010","011101101111","011101101100",
"011101101000","011101100101","011101100010","011101011111","011101011100","011101011001","011101010110","011101010010",
"011101001111","011101001100","011101001001","011101000110","011101000011","011101000000","011100111101","011100111001",
"011100110110","011100110011","011100110000","011100101101","011100101010","011100100111","011100100100","011100100000",
"011100011101","011100011010","011100010111","011100010100","011100010001","011100001110","011100001011","011100000111",
"011100000100","011100000001","011011111110","011011111011","011011111000","011011110101","011011110010","011011101111",
"011011101011","011011101000","011011100101","011011100010","011011011111","011011011100","011011011001","011011010110",
"011011010011","011011001111","011011001100","011011001001","011011000110","011011000011","011011000000","011010111101",
"011010111010","011010110111","011010110100","011010110000","011010101101","011010101010","011010100111","011010100100",
"011010100001","011010011110","011010011011","011010011000","011010010101","011010010001","011010001110","011010001011",
"011010001000","011010000101","011010000010","011001111111","011001111100","011001111001","011001110110","011001110011",
"011001110000","011001101100","011001101001","011001100110","011001100011","011001100000","011001011101","011001011010",
"011001010111","011001010100","011001010001","011001001110","011001001011","011001001000","011001000101","011001000001",
"011000111110","011000111011","011000111000","011000110101","011000110010","011000101111","011000101100","011000101001",
"011000100110","011000100011","011000100000","011000011101","011000011010","011000010111","011000010100","011000010001",
"011000001101","011000001010","011000000111","011000000100","011000000001","010111111110","010111111011","010111111000",
"010111110101","010111110010","010111101111","010111101100","010111101001","010111100110","010111100011","010111100000",
"010111011101","010111011010","010111010111","010111010100","010111010001","010111001110","010111001011","010111001000",
"010111000101","010111000010","010110111111","010110111100","010110111001","010110110110","010110110011","010110110000",
"010110101101","010110101010","010110100111","010110100100","010110100001","010110011110","010110011011","010110011000",
"010110010101","010110010010","010110001111","010110001100","010110001001","010110000110","010110000011","010110000000",
"010101111101","010101111010","010101110111","010101110100","010101110001","010101101110","010101101011","010101101000",
"010101100101","010101100010","010101011111","010101011100","010101011001","010101010110","010101010011","010101010000",
"010101001101","010101001010","010101000111","010101000100","010101000001","010100111110","010100111100","010100111001",
"010100110110","010100110011","010100110000","010100101101","010100101010","010100100111","010100100100","010100100001",
"010100011110","010100011011","010100011000","010100010101","010100010010","010100001111","010100001101","010100001010",
"010100000111","010100000100","010100000001","010011111110","010011111011","010011111000","010011110101","010011110010",
"010011101111","010011101101","010011101010","010011100111","010011100100","010011100001","010011011110","010011011011",
"010011011000","010011010101","010011010011","010011010000","010011001101","010011001010","010011000111","010011000100",
"010011000001","010010111110","010010111100","010010111001","010010110110","010010110011","010010110000","010010101101",
"010010101010","010010101000","010010100101","010010100010","010010011111","010010011100","010010011001","010010010110",
"010010010100","010010010001","010010001110","010010001011","010010001000","010010000101","010010000011","010010000000",
"010001111101","010001111010","010001110111","010001110100","010001110010","010001101111","010001101100","010001101001",
"010001100110","010001100100","010001100001","010001011110","010001011011","010001011000","010001010110","010001010011",
"010001010000","010001001101","010001001010","010001001000","010001000101","010001000010","010000111111","010000111101",
"010000111010","010000110111","010000110100","010000110010","010000101111","010000101100","010000101001","010000100110",
"010000100100","010000100001","010000011110","010000011011","010000011001","010000010110","010000010011","010000010001",
"010000001110","010000001011","010000001000","010000000110","010000000011","010000000000","001111111101","001111111011",
"001111111000","001111110101","001111110011","001111110000","001111101101","001111101010","001111101000","001111100101",
"001111100010","001111100000","001111011101","001111011010","001111011000","001111010101","001111010010","001111010000",
"001111001101","001111001010","001111001000","001111000101","001111000010","001111000000","001110111101","001110111010",
"001110111000","001110110101","001110110010","001110110000","001110101101","001110101010","001110101000","001110100101",
"001110100010","001110100000","001110011101","001110011011","001110011000","001110010101","001110010011","001110010000",
"001110001101","001110001011","001110001000","001110000110","001110000011","001110000000","001101111110","001101111011",
"001101111001","001101110110","001101110011","001101110001","001101101110","001101101100","001101101001","001101100111",
"001101100100","001101100001","001101011111","001101011100","001101011010","001101010111","001101010101","001101010010",
"001101010000","001101001101","001101001010","001101001000","001101000101","001101000011","001101000000","001100111110",
"001100111011","001100111001","001100110110","001100110100","001100110001","001100101111","001100101100","001100101010",
"001100100111","001100100101","001100100010","001100100000","001100011101","001100011011","001100011000","001100010110",
"001100010011","001100010001","001100001110","001100001100","001100001001","001100000111","001100000101","001100000010",
"001100000000","001011111101","001011111011","001011111000","001011110110","001011110011","001011110001","001011101111",
"001011101100","001011101010","001011100111","001011100101","001011100010","001011100000","001011011110","001011011011",
"001011011001","001011010110","001011010100","001011010010","001011001111","001011001101","001011001010","001011001000",
"001011000110","001011000011","001011000001","001010111111","001010111100","001010111010","001010110111","001010110101",
"001010110011","001010110000","001010101110","001010101100","001010101001","001010100111","001010100101","001010100010",
"001010100000","001010011110","001010011011","001010011001","001010010111","001010010100","001010010010","001010010000",
"001010001101","001010001011","001010001001","001010000111","001010000100","001010000010","001010000000","001001111101",
"001001111011","001001111001","001001110111","001001110100","001001110010","001001110000","001001101110","001001101011",
"001001101001","001001100111","001001100101","001001100010","001001100000","001001011110","001001011100","001001011001",
"001001010111","001001010101","001001010011","001001010001","001001001110","001001001100","001001001010","001001001000",
"001001000110","001001000011","001001000001","001000111111","001000111101","001000111011","001000111000","001000110110",
"001000110100","001000110010","001000110000","001000101110","001000101011","001000101001","001000100111","001000100101",
"001000100011","001000100001","001000011111","001000011100","001000011010","001000011000","001000010110","001000010100",
"001000010010","001000010000","001000001110","001000001100","001000001001","001000000111","001000000101","001000000011",
"001000000001","000111111111","000111111101","000111111011","000111111001","000111110111","000111110101","000111110011",
"000111110001","000111101111","000111101101","000111101010","000111101000","000111100110","000111100100","000111100010",
"000111100000","000111011110","000111011100","000111011010","000111011000","000111010110","000111010100","000111010010",
"000111010000","000111001110","000111001100","000111001010","000111001000","000111000110","000111000100","000111000010",
"000111000000","000110111110","000110111101","000110111011","000110111001","000110110111","000110110101","000110110011",
"000110110001","000110101111","000110101101","000110101011","000110101001","000110100111","000110100101","000110100011",
"000110100010","000110100000","000110011110","000110011100","000110011010","000110011000","000110010110","000110010100",
"000110010010","000110010001","000110001111","000110001101","000110001011","000110001001","000110000111","000110000101",
"000110000100","000110000010","000110000000","000101111110","000101111100","000101111010","000101111001","000101110111",
"000101110101","000101110011","000101110001","000101110000","000101101110","000101101100","000101101010","000101101000",
"000101100111","000101100101","000101100011","000101100001","000101100000","000101011110","000101011100","000101011010",
"000101011001","000101010111","000101010101","000101010011","000101010010","000101010000","000101001110","000101001100",
"000101001011","000101001001","000101000111","000101000110","000101000100","000101000010","000101000001","000100111111",
"000100111101","000100111011","000100111010","000100111000","000100110110","000100110101","000100110011","000100110001",
"000100110000","000100101110","000100101101","000100101011","000100101001","000100101000","000100100110","000100100100",
"000100100011","000100100001","000100100000","000100011110","000100011100","000100011011","000100011001","000100011000",
"000100010110","000100010100","000100010011","000100010001","000100010000","000100001110","000100001101","000100001011",
"000100001001","000100001000","000100000110","000100000101","000100000011","000100000010","000100000000","000011111111",
"000011111101","000011111100","000011111010","000011111001","000011110111","000011110110","000011110100","000011110011",
"000011110001","000011110000","000011101110","000011101101","000011101011","000011101010","000011101000","000011100111",
"000011100110","000011100100","000011100011","000011100001","000011100000","000011011110","000011011101","000011011100",
"000011011010","000011011001","000011010111","000011010110","000011010101","000011010011","000011010010","000011010000",
"000011001111","000011001110","000011001100","000011001011","000011001001","000011001000","000011000111","000011000101",
"000011000100","000011000011","000011000001","000011000000","000010111111","000010111101","000010111100","000010111011",
"000010111001","000010111000","000010110111","000010110110","000010110100","000010110011","000010110010","000010110000",
"000010101111","000010101110","000010101101","000010101011","000010101010","000010101001","000010101000","000010100110",
"000010100101","000010100100","000010100011","000010100001","000010100000","000010011111","000010011110","000010011101",
"000010011011","000010011010","000010011001","000010011000","000010010111","000010010101","000010010100","000010010011",
"000010010010","000010010001","000010010000","000010001110","000010001101","000010001100","000010001011","000010001010",
"000010001001","000010001000","000010000110","000010000101","000010000100","000010000011","000010000010","000010000001",
"000010000000","000001111111","000001111110","000001111101","000001111011","000001111010","000001111001","000001111000",
"000001110111","000001110110","000001110101","000001110100","000001110011","000001110010","000001110001","000001110000",
"000001101111","000001101110","000001101101","000001101100","000001101011","000001101010","000001101001","000001101000",
"000001100111","000001100110","000001100101","000001100100","000001100011","000001100010","000001100001","000001100000",
"000001011111","000001011110","000001011101","000001011100","000001011011","000001011010","000001011001","000001011001",
"000001011000","000001010111","000001010110","000001010101","000001010100","000001010011","000001010010","000001010001",
"000001010001","000001010000","000001001111","000001001110","000001001101","000001001100","000001001011","000001001011",
"000001001010","000001001001","000001001000","000001000111","000001000110","000001000110","000001000101","000001000100",
"000001000011","000001000010","000001000010","000001000001","000001000000","000000111111","000000111110","000000111110",
"000000111101","000000111100","000000111011","000000111011","000000111010","000000111001","000000111000","000000111000",
"000000110111","000000110110","000000110101","000000110101","000000110100","000000110011","000000110011","000000110010",
"000000110001","000000110001","000000110000","000000101111","000000101111","000000101110","000000101101","000000101101",
"000000101100","000000101011","000000101011","000000101010","000000101001","000000101001","000000101000","000000100111",
"000000100111","000000100110","000000100110","000000100101","000000100100","000000100100","000000100011","000000100011",
"000000100010","000000100010","000000100001","000000100000","000000100000","000000011111","000000011111","000000011110",
"000000011110","000000011101","000000011101","000000011100","000000011100","000000011011","000000011011","000000011010",
"000000011010","000000011001","000000011001","000000011000","000000011000","000000010111","000000010111","000000010110",
"000000010110","000000010101","000000010101","000000010100","000000010100","000000010011","000000010011","000000010011",
"000000010010","000000010010","000000010001","000000010001","000000010000","000000010000","000000010000","000000001111",
"000000001111","000000001111","000000001110","000000001110","000000001101","000000001101","000000001101","000000001100",
"000000001100","000000001100","000000001011","000000001011","000000001011","000000001010","000000001010","000000001010",
"000000001001","000000001001","000000001001","000000001000","000000001000","000000001000","000000001000","000000000111",
"000000000111","000000000111","000000000111","000000000110","000000000110","000000000110","000000000110","000000000101",
"000000000101","000000000101","000000000101","000000000100","000000000100","000000000100","000000000100","000000000100",
"000000000011","000000000011","000000000011","000000000011","000000000011","000000000010","000000000010","000000000010",
"000000000010","000000000010","000000000010","000000000010","000000000001","000000000001","000000000001","000000000001",
"000000000001","000000000001","000000000001","000000000001","000000000000","000000000000","000000000000","000000000000",
"000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000",
"000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000",
"000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000",
"000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000",
"000000000000","000000000000","000000000000","000000000000","000000000000","000000000001","000000000001","000000000001",
"000000000001","000000000001","000000000001","000000000001","000000000001","000000000010","000000000010","000000000010",
"000000000010","000000000010","000000000010","000000000010","000000000011","000000000011","000000000011","000000000011",
"000000000011","000000000100","000000000100","000000000100","000000000100","000000000100","000000000101","000000000101",
"000000000101","000000000101","000000000110","000000000110","000000000110","000000000110","000000000111","000000000111",
"000000000111","000000000111","000000001000","000000001000","000000001000","000000001000","000000001001","000000001001",
"000000001001","000000001010","000000001010","000000001010","000000001011","000000001011","000000001011","000000001100",
"000000001100","000000001100","000000001101","000000001101","000000001101","000000001110","000000001110","000000001111",
"000000001111","000000001111","000000010000","000000010000","000000010000","000000010001","000000010001","000000010010",
"000000010010","000000010011","000000010011","000000010011","000000010100","000000010100","000000010101","000000010101",
"000000010110","000000010110","000000010111","000000010111","000000011000","000000011000","000000011001","000000011001",
"000000011010","000000011010","000000011011","000000011011","000000011100","000000011100","000000011101","000000011101",
"000000011110","000000011110","000000011111","000000011111","000000100000","000000100000","000000100001","000000100010",
"000000100010","000000100011","000000100011","000000100100","000000100100","000000100101","000000100110","000000100110",
"000000100111","000000100111","000000101000","000000101001","000000101001","000000101010","000000101011","000000101011",
"000000101100","000000101101","000000101101","000000101110","000000101111","000000101111","000000110000","000000110001",
"000000110001","000000110010","000000110011","000000110011","000000110100","000000110101","000000110101","000000110110",
"000000110111","000000111000","000000111000","000000111001","000000111010","000000111011","000000111011","000000111100",
"000000111101","000000111110","000000111110","000000111111","000001000000","000001000001","000001000010","000001000010",
"000001000011","000001000100","000001000101","000001000110","000001000110","000001000111","000001001000","000001001001",
"000001001010","000001001011","000001001011","000001001100","000001001101","000001001110","000001001111","000001010000",
"000001010001","000001010001","000001010010","000001010011","000001010100","000001010101","000001010110","000001010111",
"000001011000","000001011001","000001011001","000001011010","000001011011","000001011100","000001011101","000001011110",
"000001011111","000001100000","000001100001","000001100010","000001100011","000001100100","000001100101","000001100110",
"000001100111","000001101000","000001101001","000001101010","000001101011","000001101100","000001101101","000001101110",
"000001101111","000001110000","000001110001","000001110010","000001110011","000001110100","000001110101","000001110110",
"000001110111","000001111000","000001111001","000001111010","000001111011","000001111101","000001111110","000001111111",
"000010000000","000010000001","000010000010","000010000011","000010000100","000010000101","000010000110","000010001000",
"000010001001","000010001010","000010001011","000010001100","000010001101","000010001110","000010010000","000010010001",
"000010010010","000010010011","000010010100","000010010101","000010010111","000010011000","000010011001","000010011010",
"000010011011","000010011101","000010011110","000010011111","000010100000","000010100001","000010100011","000010100100",
"000010100101","000010100110","000010101000","000010101001","000010101010","000010101011","000010101101","000010101110",
"000010101111","000010110000","000010110010","000010110011","000010110100","000010110110","000010110111","000010111000",
"000010111001","000010111011","000010111100","000010111101","000010111111","000011000000","000011000001","000011000011",
"000011000100","000011000101","000011000111","000011001000","000011001001","000011001011","000011001100","000011001110",
"000011001111","000011010000","000011010010","000011010011","000011010101","000011010110","000011010111","000011011001",
"000011011010","000011011100","000011011101","000011011110","000011100000","000011100001","000011100011","000011100100",
"000011100110","000011100111","000011101000","000011101010","000011101011","000011101101","000011101110","000011110000",
"000011110001","000011110011","000011110100","000011110110","000011110111","000011111001","000011111010","000011111100",
"000011111101","000011111111","000100000000","000100000010","000100000011","000100000101","000100000110","000100001000",
"000100001001","000100001011","000100001101","000100001110","000100010000","000100010001","000100010011","000100010100",
"000100010110","000100011000","000100011001","000100011011","000100011100","000100011110","000100100000","000100100001",
"000100100011","000100100100","000100100110","000100101000","000100101001","000100101011","000100101101","000100101110",
"000100110000","000100110001","000100110011","000100110101","000100110110","000100111000","000100111010","000100111011",
"000100111101","000100111111","000101000001","000101000010","000101000100","000101000110","000101000111","000101001001",
"000101001011","000101001100","000101001110","000101010000","000101010010","000101010011","000101010101","000101010111",
"000101011001","000101011010","000101011100","000101011110","000101100000","000101100001","000101100011","000101100101",
"000101100111","000101101000","000101101010","000101101100","000101101110","000101110000","000101110001","000101110011",
"000101110101","000101110111","000101111001","000101111010","000101111100","000101111110","000110000000","000110000010",
"000110000100","000110000101","000110000111","000110001001","000110001011","000110001101","000110001111","000110010001",
"000110010010","000110010100","000110010110","000110011000","000110011010","000110011100","000110011110","000110100000",
"000110100010","000110100011","000110100101","000110100111","000110101001","000110101011","000110101101","000110101111",
"000110110001","000110110011","000110110101","000110110111","000110111001","000110111011","000110111101","000110111110",
"000111000000","000111000010","000111000100","000111000110","000111001000","000111001010","000111001100","000111001110",
"000111010000","000111010010","000111010100","000111010110","000111011000","000111011010","000111011100","000111011110",
"000111100000","000111100010","000111100100","000111100110","000111101000","000111101010","000111101101","000111101111",
"000111110001","000111110011","000111110101","000111110111","000111111001","000111111011","000111111101","000111111111",
"001000000001","001000000011","001000000101","001000000111","001000001001","001000001100","001000001110","001000010000",
"001000010010","001000010100","001000010110","001000011000","001000011010","001000011100","001000011111","001000100001",
"001000100011","001000100101","001000100111","001000101001","001000101011","001000101110","001000110000","001000110010",
"001000110100","001000110110","001000111000","001000111011","001000111101","001000111111","001001000001","001001000011",
"001001000110","001001001000","001001001010","001001001100","001001001110","001001010001","001001010011","001001010101",
"001001010111","001001011001","001001011100","001001011110","001001100000","001001100010","001001100101","001001100111",
"001001101001","001001101011","001001101110","001001110000","001001110010","001001110100","001001110111","001001111001",
"001001111011","001001111101","001010000000","001010000010","001010000100","001010000111","001010001001","001010001011",
"001010001101","001010010000","001010010010","001010010100","001010010111","001010011001","001010011011","001010011110",
"001010100000","001010100010","001010100101","001010100111","001010101001","001010101100","001010101110","001010110000",
"001010110011","001010110101","001010110111","001010111010","001010111100","001010111111","001011000001","001011000011",
"001011000110","001011001000","001011001010","001011001101","001011001111","001011010010","001011010100","001011010110",
"001011011001","001011011011","001011011110","001011100000","001011100010","001011100101","001011100111","001011101010",
"001011101100","001011101111","001011110001","001011110011","001011110110","001011111000","001011111011","001011111101",
"001100000000","001100000010","001100000101","001100000111","001100001001","001100001100","001100001110","001100010001",
"001100010011","001100010110","001100011000","001100011011","001100011101","001100100000","001100100010","001100100101",
"001100100111","001100101010","001100101100","001100101111","001100110001","001100110100","001100110110","001100111001",
"001100111011","001100111110","001101000000","001101000011","001101000101","001101001000","001101001010","001101001101",
"001101010000","001101010010","001101010101","001101010111","001101011010","001101011100","001101011111","001101100001",
"001101100100","001101100111","001101101001","001101101100","001101101110","001101110001","001101110011","001101110110",
"001101111001","001101111011","001101111110","001110000000","001110000011","001110000110","001110001000","001110001011",
"001110001101","001110010000","001110010011","001110010101","001110011000","001110011011","001110011101","001110100000",
"001110100010","001110100101","001110101000","001110101010","001110101101","001110110000","001110110010","001110110101",
"001110111000","001110111010","001110111101","001111000000","001111000010","001111000101","001111001000","001111001010",
"001111001101","001111010000","001111010010","001111010101","001111011000","001111011010","001111011101","001111100000",
"001111100010","001111100101","001111101000","001111101010","001111101101","001111110000","001111110011","001111110101",
"001111111000","001111111011","001111111101","010000000000","010000000011","010000000110","010000001000","010000001011",
"010000001110","010000010001","010000010011","010000010110","010000011001","010000011011","010000011110","010000100001",
"010000100100","010000100110","010000101001","010000101100","010000101111","010000110010","010000110100","010000110111",
"010000111010","010000111101","010000111111","010001000010","010001000101","010001001000","010001001010","010001001101",
"010001010000","010001010011","010001010110","010001011000","010001011011","010001011110","010001100001","010001100100",
"010001100110","010001101001","010001101100","010001101111","010001110010","010001110100","010001110111","010001111010",
"010001111101","010010000000","010010000011","010010000101","010010001000","010010001011","010010001110","010010010001",
"010010010100","010010010110","010010011001","010010011100","010010011111","010010100010","010010100101","010010101000",
"010010101010","010010101101","010010110000","010010110011","010010110110","010010111001","010010111100","010010111110",
"010011000001","010011000100","010011000111","010011001010","010011001101","010011010000","010011010011","010011010101",
"010011011000","010011011011","010011011110","010011100001","010011100100","010011100111","010011101010","010011101101",
"010011101111","010011110010","010011110101","010011111000","010011111011","010011111110","010100000001","010100000100",
"010100000111","010100001010","010100001101","010100001111","010100010010","010100010101","010100011000","010100011011",
"010100011110","010100100001","010100100100","010100100111","010100101010","010100101101","010100110000","010100110011",
"010100110110","010100111001","010100111100","010100111110","010101000001","010101000100","010101000111","010101001010",
"010101001101","010101010000","010101010011","010101010110","010101011001","010101011100","010101011111","010101100010",
"010101100101","010101101000","010101101011","010101101110","010101110001","010101110100","010101110111","010101111010",
"010101111101","010110000000","010110000011","010110000110","010110001001","010110001100","010110001111","010110010010",
"010110010101","010110011000","010110011011","010110011110","010110100001","010110100100","010110100111","010110101010",
"010110101101","010110110000","010110110011","010110110110","010110111001","010110111100","010110111111","010111000010",
"010111000101","010111001000","010111001011","010111001110","010111010001","010111010100","010111010111","010111011010",
"010111011101","010111100000","010111100011","010111100110","010111101001","010111101100","010111101111","010111110010",
"010111110101","010111111000","010111111011","010111111110","011000000001","011000000100","011000000111","011000001010",
"011000001101","011000010001","011000010100","011000010111","011000011010","011000011101","011000100000","011000100011",
"011000100110","011000101001","011000101100","011000101111","011000110010","011000110101","011000111000","011000111011",
"011000111110","011001000001","011001000101","011001001000","011001001011","011001001110","011001010001","011001010100",
"011001010111","011001011010","011001011101","011001100000","011001100011","011001100110","011001101001","011001101100",
"011001110000","011001110011","011001110110","011001111001","011001111100","011001111111","011010000010","011010000101",
"011010001000","011010001011","011010001110","011010010001","011010010101","011010011000","011010011011","011010011110",
"011010100001","011010100100","011010100111","011010101010","011010101101","011010110000","011010110100","011010110111",
"011010111010","011010111101","011011000000","011011000011","011011000110","011011001001","011011001100","011011001111",
"011011010011","011011010110","011011011001","011011011100","011011011111","011011100010","011011100101","011011101000",
"011011101011","011011101111","011011110010","011011110101","011011111000","011011111011","011011111110","011100000001",
"011100000100","011100000111","011100001011","011100001110","011100010001","011100010100","011100010111","011100011010",
"011100011101","011100100000","011100100100","011100100111","011100101010","011100101101","011100110000","011100110011",
"011100110110","011100111001","011100111101","011101000000","011101000011","011101000110","011101001001","011101001100",
"011101001111","011101010010","011101010110","011101011001","011101011100","011101011111","011101100010","011101100101",
"011101101000","011101101100","011101101111","011101110010","011101110101","011101111000","011101111011","011101111110",
"011110000001","011110000101","011110001000","011110001011","011110001110","011110010001","011110010100","011110010111",
"011110011011","011110011110","011110100001","011110100100","011110100111","011110101010","011110101101","011110110000",
"011110110100","011110110111","011110111010","011110111101","011111000000","011111000011","011111000110","011111001010",
"011111001101","011111010000","011111010011","011111010110","011111011001","011111011100","011111100000","011111100011",
"011111100110","011111101001","011111101100","011111101111","011111110010","011111110110","011111111001","011111111100"
);

-- LUT index and sine value
signal lut_index : integer range 0 to 4095; -- 12-bit range
signal sine_value: STD_LOGIC_VECTOR(11 downto 0);

-- Horizontal and Vertical counters
signal h_counter : integer range 0 to HOR_RES + HOR_FRONT + HOR_SYNC + HOR_BACK := 0;
signal v_counter : integer range 0 to VER_RES + VER_FRONT + VER_SYNC + VER_BACK := 0;

-- Pixel valid signal
signal pixel_valid : std_logic;

-- Compute LUT indices based on h_counter for different colors
signal lut_index_r : integer range 0 to 4095; -- 12-bit range
signal lut_index_g : integer range 0 to 4095; -- 12-bit range
signal lut_index_b : integer range 0 to 4095; -- 12-bit range

signal sine_value_r: STD_LOGIC_VECTOR(11 downto 0);
signal sine_value_g: STD_LOGIC_VECTOR(11 downto 0);
signal sine_value_b: STD_LOGIC_VECTOR(11 downto 0);

begin

-- Compute LUT indices with different phase offsets
lut_index_r <= (h_counter * 4096) / HOR_RES;
lut_index_g <= (lut_index_r + 1365) mod 4096; -- Offset by 1/3 of the wave
lut_index_b <= (lut_index_r + 2730) mod 4096; -- Offset by 2/3 of the wave


-- Get sine values from LUT
sine_value_r <= SIN_LUT(lut_index_r);
sine_value_g <= SIN_LUT(lut_index_g);
sine_value_b <= SIN_LUT(lut_index_b);


-- Horizontal Counter
H_COUNT: process(clock_50, reset)
begin
  if reset = '1' then
    h_counter <= 0;
  elsif rising_edge(clock_50) then
    if h_counter = HOR_RES + HOR_FRONT + HOR_SYNC + HOR_BACK - 1 then
      h_counter <= 0;
    else
      h_counter <= h_counter + 1;
    end if;
  end if;
end process H_COUNT;

-- Vertical Counter
V_COUNT: process(clock_50, reset)
begin
  if reset = '1' then
    v_counter <= 0;
  elsif rising_edge(clock_50) then
    if h_counter = HOR_RES + HOR_FRONT + HOR_SYNC + HOR_BACK - 1 then
      if v_counter = VER_RES + VER_FRONT + VER_SYNC + VER_BACK - 1 then
        v_counter <= 0;
      else
        v_counter <= v_counter + 1;
      end if;
    end if;
  end if;
end process V_COUNT;

-- Generate sync signals
vga_hs <= '1' when h_counter < HOR_RES + HOR_FRONT or h_counter >= HOR_RES + HOR_FRONT + HOR_SYNC else '0';
vga_vs <= '1' when v_counter < VER_RES + VER_FRONT or v_counter >= VER_RES + VER_FRONT + VER_SYNC else '0';

-- Generate pixel_valid signal
pixel_valid <= '1' when h_counter < HOR_RES and v_counter < VER_RES else '0';

-- Add a process to handle the color outputs based on the state
process(clock_50, reset)
begin
    if reset = '1' then
        vga_r <= (others => '0');
        vga_g <= (others => '0');
        vga_b <= (others => '0');
    elsif rising_edge(clock_50) then
        if current_state = ready then
            -- Output rainbow colors
            if pixel_valid = '1' then
                vga_r <= sine_value_r;
                vga_g <= sine_value_g;
                vga_b <= sine_value_b;
            else
                vga_r <= (others => '0');
                vga_g <= (others => '0');
                vga_b <= (others => '0');
            end if;
        elsif current_state = fail then
            -- Output solid red color
            if pixel_valid = '1' then
                vga_r <= "111111111111";
            else
                vga_r <= (others => '0');
            end if;
            vga_g <= (others => '0');
            vga_b <= (others => '0');
			elsif current_state = yes then
            -- Output solid green color
            if pixel_valid = '1' then
                vga_g <= "111111111111";
            else
                vga_g <= (others => '0');
            end if;
            vga_r <= (others => '0');
            vga_b <= (others => '0');
        else
            -- Default behavior
            vga_r <= "000000000000";
            vga_b <= "111111111111";
            vga_g <= "111111111111";
        end if;
    end if;
end process;

end Behavioral;

